`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    17:20:06 10/22/2016
// Design Name:
// Module Name:    Top_Module
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module Top_Module(RST,PC_LIMIT,CLK,
EX_FLAG,
LED_STATUS,
REGISTER_A,REGISTER_B,
PC_COUNTER);

output LED_STATUS;
wire [16:0]temp_alu_result;
wire carry,zero;
input RST;
input[2:0]PC_LIMIT;
input CLK;
wire IFF;

wire [1:0]SELECT;
wire SELECT_DEMUX;
wire [1:0] SELECT2;
wire DECODE_FLAG;

wire [15:0] DATA_IN;
wire WRITE_ENABLE;
wire REG_WRITE_ENABLE;
wire DATA_WRITE_ENABLE;

wire [11:0] PC_ADDRESS;
wire [15:0] DATA_REGISTER_SET;
wire [15:0] ALU_RESULT_OUT;

wire [7:0] ALU_OPCODE2;
wire [11:0] ADDRESS;
wire [15:0] DATA_OUT;
wire [2:0] OPERAND1;
wire [2:0] OPERAND2;
wire [2:0] DESTINATION;
wire [11:0] DATA_ADDR;
wire [15:0] WRITE_DATA;
wire [15:0] READ_A;
wire [15:0] READ_B;
wire [7:0] OPCODE2;

wire [11:0] ADDR;
wire [3:0] OPCODE1;

inout EX_FLAG;
//wire EX_FLAG;
wire [15:0] DATA_M_OUT;
wire [15:0] DATA_INPUT;
wire [15:0] REG_DATA_OUT;

wire STACK_EN;
wire [15:0] STACK_IN;
wire [11:0] SP_OUT;

wire [1:0] JMP_EN;
wire [11:0] JMP_ADDR;

wire [1:0] STACK_MUX_SEL;
wire [15:0] STACK_REG;

wire STACK_PC_EN;
wire [15:0] DEMUX_PC_IN;
wire [15:0] REG_MUX_IN;

wire [15:0] ZERO_CARRY_IEN;
wire ZC_FLAG;
wire [2:0] INTERRUPT_COUNTER;
output [15:0]REGISTER_A;
output [15:0]REGISTER_B;

//wire [15:0]REGISTER_A;
//wire [15:0]REGISTER_B;

wire [15:0]REGISTER_C;
wire [15:0]REGISTER_Z;
inout [4:0]PC_COUNTER;
wire RET_FLAG;

A5_PC_BLOCK uut1(PC_COUNTER,REGISTER_A,REGISTER_C,REGISTER_Z,LED_STATUS,CLK,RST,PC_LIMIT,EX_FLAG,RET_FLAG,PC_ADDRESS,JMP_EN,JMP_ADDR,DEMUX_PC_IN,
ZC_FLAG,IFF,INTERRUPT_COUNTER);
A5_memory uut2(DATA_IN,WRITE_ENABLE,PC_ADDRESS,CLK,DATA_OUT);//MEM);
A5_INST_DECODE uut3(ZERO_CARRY_IEN,DATA_OUT,CLK,OPERAND1,OPERAND2,DESTINATION,DATA_ADDR,OPCODE2,DECODE_FLAG,
SELECT,SELECT2,SELECT_DEMUX,ADDR,OPCODE1,JMP_ADDR, STACK_MUX_SEL,STACK_PC_EN,ZC_FLAG, IFF, INTERRUPT_COUNTER, EX_FLAG);
A5_register_set uut4(REGISTER_A,REGISTER_B,REGISTER_C,REGISTER_Z,CLK,OPERAND1,OPERAND2,DESTINATION,WRITE_DATA,REG_WRITE_ENABLE,REG_DATA_OUT,READ_B,DATA_REGISTER_SET,ZERO_CARRY_IEN,temp_alu_result);
A5_Data_Memory uut5(DATA_INPUT, DATA_WRITE_ENABLE, ADDRESS, CLK, DATA_M_OUT);//,DATA_MEM);
A5_ALU uut6(CLK,READ_A,READ_B, ALU_OPCODE2,ALU_RESULT_OUT,carry,zero,temp_alu_result);
ALU_DATA_MEM_MUX uut7(CLK,SELECT, DATA_M_OUT,ALU_RESULT_OUT,WRITE_DATA, REG_MUX_IN);
A5_DATA_ALU_DEMUX uu8(CLK, DATA_ADDR, OPCODE2, SELECT_DEMUX, ADDRESS, ALU_OPCODE2 );
A5_CONTROL_UNIT uut9(REGISTER_C,REGISTER_Z,PC_COUNTER,RST, CLK, DECODE_FLAG,REG_WRITE_ENABLE, EX_FLAG,RET_FLAG,ADDR,OPCODE1,DATA_WRITE_ENABLE,OPCODE2, STACK_EN,JMP_EN, IFF, INTERRUPT_COUNTER);
A5_DATA_ALU_REG_DEMUX uut10(CLK, REG_DATA_OUT, SELECT2, DATA_INPUT, READ_A, STACK_REG);
A5_STACK uut11(CLK,STACK_IN,REG_MUX_IN,STACK_EN,SP_OUT,STACK_PC_EN, DEMUX_PC_IN);
A5_STACK_MUX uut12(CLK, PC_ADDRESS, STACK_REG, STACK_IN, STACK_MUX_SEL);

endmodule
